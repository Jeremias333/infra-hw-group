module mult #(parameter N=2)
	(input start, rst, 
	output reg [7:0] saida);

	while(incrementar <= b) begin
		saida += a;
		incrementar++;
	end

endmodule
