/*
-Nome do grupo: LearnWARE 
-Questão de número: 4
-Data: 27/05/2022
-Atividade de número: 3
-Disciplina: Infraestrutura de Hardware
-Professor: Vitor Coutinho
-Semestre Letivo: 3º semestre
-Turma: B
-Alunos: Paulo Guerreiro, Elder Lamarck, Jacquelin Busch, Jeremias Oliveira
-Objetivo do algoritmo: É uma multiplicar sem usar o operador de multiplicação em verilog.
*/
module mult #(parameter N=2)
	(input start, rst, 
	output reg [7:0] saida);

	while(incrementar <= b) begin
		saida += a;
		incrementar++;
	end

endmodule
